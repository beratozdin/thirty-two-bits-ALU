`define DELAY 20
module thirty_two_alu_testbench(); 
reg [31:0] Ai;
reg [31:0] Bi;
reg Op2,Op1,Op0;
wire [31:0] Ri;
wire Cout,Vout,Z;

thirty_two_alu gate_thirty_alu(Ai,Bi,Ri,Cout,Vout,Z,Op2,Op1,Op0);

initial begin
Ai=32'b01101111000011110000111101011010; Bi=32'b01101111000011110000111101011010; Op2=1'b0; Op1=1'b0; Op0=1'b0;
#`DELAY;
Ai=32'b01101111000011110000111101011010; Bi=32'b01101111000011110000111101011010; Op2=1'b0; Op1=1'b0; Op0=1'b1;
#`DELAY;
Ai=32'b01101111000011110000111101011010; Bi=32'b01101111000011110000111101011010; Op2=1'b0; Op1=1'b1; Op0=1'b0;
#`DELAY;
Ai=32'b01101111000011110000111101011010; Bi=32'b01101111000011110000111101011010; Op2=1'b1; Op1=1'b1; Op0=1'b0;
#`DELAY;
Ai=32'b01101111000011110000111101011010; Bi=32'b01101111000011110000111101011010; Op2=1'b1; Op1=1'b1; Op0=1'b1;

#`DELAY;
Ai=32'b11101111000010110100110101011010; Bi=32'b01101111010011110000101101011010; Op2=1'b0; Op1=1'b0; Op0=1'b0;
#`DELAY;
Ai=32'b11101111000010110100110101011010; Bi=32'b01101111010011110000101101011010; Op2=1'b0; Op1=1'b0; Op0=1'b1;
#`DELAY;
Ai=32'b11101111000010110100110101011010; Bi=32'b01101111010011110000101101011010; Op2=1'b0; Op1=1'b1; Op0=1'b0;
#`DELAY;
Ai=32'b11101111000010110100110101011010; Bi=32'b01101111010011110000101101011010; Op2=1'b1; Op1=1'b1; Op0=1'b0;
#`DELAY;
Ai=32'b11101111000010110100110101011010; Bi=32'b01101111010011110000101101011010; Op2=1'b1; Op1=1'b1; Op0=1'b1;

#`DELAY;
Ai=32'b01101111000010110110111101011010; Bi=32'b01101011000011110000111101011010; Op2=1'b0; Op1=1'b0; Op0=1'b0;
#`DELAY;
Ai=32'b01101111000010110110111101011010; Bi=32'b01101011000011110000111101011010; Op2=1'b0; Op1=1'b0; Op0=1'b1;
#`DELAY;
Ai=32'b01101111000010110110111101011010; Bi=32'b01101011000011110000111101011010; Op2=1'b0; Op1=1'b1; Op0=1'b0;
#`DELAY;
Ai=32'b01101111000010110110111101011010; Bi=32'b01101011000011110000111101011010; Op2=1'b1; Op1=1'b1; Op0=1'b0;
#`DELAY;
Ai=32'b01101111000010110110111101011010; Bi=32'b01101011000011110000111101011010; Op2=1'b1; Op1=1'b1; Op0=1'b1;

end

initial
begin
$monitor("time = %2d, Ai=%32b, Bi=%32b, Ri=%32b, Op2=%1b, Op1=%1b, Op0=%1b, Cout=%1b, Vout=%1b, Z=%1b", $time, Ai, Bi, Ri, Op2, Op1, Op0,Cout,Vout,Z);
end

endmodule 